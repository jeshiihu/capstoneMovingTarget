-- soc_system.vhd

-- Generated using ACDS version 17.0 602

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_system is
	port (
		clk_clk                          : in    std_logic                     := '0';             --                       clk.clk
		easy_driver_x_conduit_end_dir    : out   std_logic;                                        -- easy_driver_x_conduit_end.dir
		easy_driver_x_conduit_end_step   : out   std_logic;                                        --                          .step
		easy_driver_x_conduit_end_enable : out   std_logic;                                        --                          .enable
		easy_driver_y_conduit_end_dir    : out   std_logic;                                        -- easy_driver_y_conduit_end.dir
		easy_driver_y_conduit_end_step   : out   std_logic;                                        --                          .step
		easy_driver_y_conduit_end_enable : out   std_logic;                                        --                          .enable
		hps_io_hps_io_emac1_inst_TX_CLK  : out   std_logic;                                        --                    hps_io.hps_io_emac1_inst_TX_CLK
		hps_io_hps_io_emac1_inst_TXD0    : out   std_logic;                                        --                          .hps_io_emac1_inst_TXD0
		hps_io_hps_io_emac1_inst_TXD1    : out   std_logic;                                        --                          .hps_io_emac1_inst_TXD1
		hps_io_hps_io_emac1_inst_TXD2    : out   std_logic;                                        --                          .hps_io_emac1_inst_TXD2
		hps_io_hps_io_emac1_inst_TXD3    : out   std_logic;                                        --                          .hps_io_emac1_inst_TXD3
		hps_io_hps_io_emac1_inst_RXD0    : in    std_logic                     := '0';             --                          .hps_io_emac1_inst_RXD0
		hps_io_hps_io_emac1_inst_MDIO    : inout std_logic                     := '0';             --                          .hps_io_emac1_inst_MDIO
		hps_io_hps_io_emac1_inst_MDC     : out   std_logic;                                        --                          .hps_io_emac1_inst_MDC
		hps_io_hps_io_emac1_inst_RX_CTL  : in    std_logic                     := '0';             --                          .hps_io_emac1_inst_RX_CTL
		hps_io_hps_io_emac1_inst_TX_CTL  : out   std_logic;                                        --                          .hps_io_emac1_inst_TX_CTL
		hps_io_hps_io_emac1_inst_RX_CLK  : in    std_logic                     := '0';             --                          .hps_io_emac1_inst_RX_CLK
		hps_io_hps_io_emac1_inst_RXD1    : in    std_logic                     := '0';             --                          .hps_io_emac1_inst_RXD1
		hps_io_hps_io_emac1_inst_RXD2    : in    std_logic                     := '0';             --                          .hps_io_emac1_inst_RXD2
		hps_io_hps_io_emac1_inst_RXD3    : in    std_logic                     := '0';             --                          .hps_io_emac1_inst_RXD3
		hps_io_hps_io_sdio_inst_CMD      : inout std_logic                     := '0';             --                          .hps_io_sdio_inst_CMD
		hps_io_hps_io_sdio_inst_D0       : inout std_logic                     := '0';             --                          .hps_io_sdio_inst_D0
		hps_io_hps_io_sdio_inst_D1       : inout std_logic                     := '0';             --                          .hps_io_sdio_inst_D1
		hps_io_hps_io_sdio_inst_CLK      : out   std_logic;                                        --                          .hps_io_sdio_inst_CLK
		hps_io_hps_io_sdio_inst_D2       : inout std_logic                     := '0';             --                          .hps_io_sdio_inst_D2
		hps_io_hps_io_sdio_inst_D3       : inout std_logic                     := '0';             --                          .hps_io_sdio_inst_D3
		hps_io_hps_io_usb1_inst_D0       : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D0
		hps_io_hps_io_usb1_inst_D1       : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D1
		hps_io_hps_io_usb1_inst_D2       : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D2
		hps_io_hps_io_usb1_inst_D3       : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D3
		hps_io_hps_io_usb1_inst_D4       : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D4
		hps_io_hps_io_usb1_inst_D5       : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D5
		hps_io_hps_io_usb1_inst_D6       : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D6
		hps_io_hps_io_usb1_inst_D7       : inout std_logic                     := '0';             --                          .hps_io_usb1_inst_D7
		hps_io_hps_io_usb1_inst_CLK      : in    std_logic                     := '0';             --                          .hps_io_usb1_inst_CLK
		hps_io_hps_io_usb1_inst_STP      : out   std_logic;                                        --                          .hps_io_usb1_inst_STP
		hps_io_hps_io_usb1_inst_DIR      : in    std_logic                     := '0';             --                          .hps_io_usb1_inst_DIR
		hps_io_hps_io_usb1_inst_NXT      : in    std_logic                     := '0';             --                          .hps_io_usb1_inst_NXT
		hps_io_hps_io_spim1_inst_CLK     : out   std_logic;                                        --                          .hps_io_spim1_inst_CLK
		hps_io_hps_io_spim1_inst_MOSI    : out   std_logic;                                        --                          .hps_io_spim1_inst_MOSI
		hps_io_hps_io_spim1_inst_MISO    : in    std_logic                     := '0';             --                          .hps_io_spim1_inst_MISO
		hps_io_hps_io_spim1_inst_SS0     : out   std_logic;                                        --                          .hps_io_spim1_inst_SS0
		hps_io_hps_io_uart0_inst_RX      : in    std_logic                     := '0';             --                          .hps_io_uart0_inst_RX
		hps_io_hps_io_uart0_inst_TX      : out   std_logic;                                        --                          .hps_io_uart0_inst_TX
		hps_io_hps_io_i2c0_inst_SDA      : inout std_logic                     := '0';             --                          .hps_io_i2c0_inst_SDA
		hps_io_hps_io_i2c0_inst_SCL      : inout std_logic                     := '0';             --                          .hps_io_i2c0_inst_SCL
		hps_io_hps_io_i2c1_inst_SDA      : inout std_logic                     := '0';             --                          .hps_io_i2c1_inst_SDA
		hps_io_hps_io_i2c1_inst_SCL      : inout std_logic                     := '0';             --                          .hps_io_i2c1_inst_SCL
		hps_io_hps_io_gpio_inst_GPIO09   : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO09
		hps_io_hps_io_gpio_inst_GPIO35   : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO35
		hps_io_hps_io_gpio_inst_GPIO40   : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO40
		hps_io_hps_io_gpio_inst_GPIO48   : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO48
		hps_io_hps_io_gpio_inst_GPIO53   : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO53
		hps_io_hps_io_gpio_inst_GPIO54   : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO54
		hps_io_hps_io_gpio_inst_GPIO61   : inout std_logic                     := '0';             --                          .hps_io_gpio_inst_GPIO61
		memory_mem_a                     : out   std_logic_vector(14 downto 0);                    --                    memory.mem_a
		memory_mem_ba                    : out   std_logic_vector(2 downto 0);                     --                          .mem_ba
		memory_mem_ck                    : out   std_logic;                                        --                          .mem_ck
		memory_mem_ck_n                  : out   std_logic;                                        --                          .mem_ck_n
		memory_mem_cke                   : out   std_logic;                                        --                          .mem_cke
		memory_mem_cs_n                  : out   std_logic;                                        --                          .mem_cs_n
		memory_mem_ras_n                 : out   std_logic;                                        --                          .mem_ras_n
		memory_mem_cas_n                 : out   std_logic;                                        --                          .mem_cas_n
		memory_mem_we_n                  : out   std_logic;                                        --                          .mem_we_n
		memory_mem_reset_n               : out   std_logic;                                        --                          .mem_reset_n
		memory_mem_dq                    : inout std_logic_vector(31 downto 0) := (others => '0'); --                          .mem_dq
		memory_mem_dqs                   : inout std_logic_vector(3 downto 0)  := (others => '0'); --                          .mem_dqs
		memory_mem_dqs_n                 : inout std_logic_vector(3 downto 0)  := (others => '0'); --                          .mem_dqs_n
		memory_mem_odt                   : out   std_logic;                                        --                          .mem_odt
		memory_mem_dm                    : out   std_logic_vector(3 downto 0);                     --                          .mem_dm
		memory_oct_rzqin                 : in    std_logic                     := '0';             --                          .oct_rzqin
		reset_reset_n                    : in    std_logic                     := '0'              --                     reset.reset_n
	);
end entity soc_system;

architecture rtl of soc_system is
	component Easy_Driver is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset_n            : in  std_logic                     := 'X';             -- reset_n
			conduit_end_dir    : out std_logic;                                        -- dir
			conduit_end_step   : out std_logic;                                        -- step
			conduit_end_enable : out std_logic;                                        -- enable
			step_read_n        : in  std_logic                     := 'X';             -- read_n
			step_readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			step_write_n       : in  std_logic                     := 'X';             -- write_n
			step_writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			dir_read_n         : in  std_logic                     := 'X';             -- read_n
			dir_readdata       : out std_logic_vector(7 downto 0);                     -- readdata
			dir_write_n        : in  std_logic                     := 'X';             -- write_n
			dir_writedata      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			period_read_n      : in  std_logic                     := 'X';             -- read_n
			period_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			period_write_n     : in  std_logic                     := 'X';             -- write_n
			period_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			duty_read_n        : in  std_logic                     := 'X';             -- read_n
			duty_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			duty_write_n       : in  std_logic                     := 'X';             -- write_n
			duty_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- writedata
		);
	end component Easy_Driver;

	component soc_system_hps_0 is
		generic (
			F2S_Width : integer := 2;
			S2F_Width : integer := 2
		);
		port (
			mem_a                    : out   std_logic_vector(14 downto 0);                    -- mem_a
			mem_ba                   : out   std_logic_vector(2 downto 0);                     -- mem_ba
			mem_ck                   : out   std_logic;                                        -- mem_ck
			mem_ck_n                 : out   std_logic;                                        -- mem_ck_n
			mem_cke                  : out   std_logic;                                        -- mem_cke
			mem_cs_n                 : out   std_logic;                                        -- mem_cs_n
			mem_ras_n                : out   std_logic;                                        -- mem_ras_n
			mem_cas_n                : out   std_logic;                                        -- mem_cas_n
			mem_we_n                 : out   std_logic;                                        -- mem_we_n
			mem_reset_n              : out   std_logic;                                        -- mem_reset_n
			mem_dq                   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			mem_odt                  : out   std_logic;                                        -- mem_odt
			mem_dm                   : out   std_logic_vector(3 downto 0);                     -- mem_dm
			oct_rzqin                : in    std_logic                     := 'X';             -- oct_rzqin
			hps_io_emac1_inst_TX_CLK : out   std_logic;                                        -- hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   : out   std_logic;                                        -- hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   : out   std_logic;                                        -- hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   : out   std_logic;                                        -- hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   : out   std_logic;                                        -- hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   : inout std_logic                     := 'X';             -- hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    : out   std_logic;                                        -- hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL : out   std_logic;                                        -- hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   : in    std_logic                     := 'X';             -- hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     : inout std_logic                     := 'X';             -- hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     : out   std_logic;                                        -- hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      : inout std_logic                     := 'X';             -- hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      : inout std_logic                     := 'X';             -- hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     : out   std_logic;                                        -- hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     : in    std_logic                     := 'X';             -- hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    : out   std_logic;                                        -- hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   : out   std_logic;                                        -- hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   : in    std_logic                     := 'X';             -- hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    : out   std_logic;                                        -- hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     : in    std_logic                     := 'X';             -- hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     : out   std_logic;                                        -- hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     : inout std_logic                     := 'X';             -- hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO48  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  : inout std_logic                     := 'X';             -- hps_io_gpio_inst_GPIO61
			h2f_rst_n                : out   std_logic;                                        -- reset_n
			h2f_lw_axi_clk           : in    std_logic                     := 'X';             -- clk
			h2f_lw_AWID              : out   std_logic_vector(11 downto 0);                    -- awid
			h2f_lw_AWADDR            : out   std_logic_vector(20 downto 0);                    -- awaddr
			h2f_lw_AWLEN             : out   std_logic_vector(3 downto 0);                     -- awlen
			h2f_lw_AWSIZE            : out   std_logic_vector(2 downto 0);                     -- awsize
			h2f_lw_AWBURST           : out   std_logic_vector(1 downto 0);                     -- awburst
			h2f_lw_AWLOCK            : out   std_logic_vector(1 downto 0);                     -- awlock
			h2f_lw_AWCACHE           : out   std_logic_vector(3 downto 0);                     -- awcache
			h2f_lw_AWPROT            : out   std_logic_vector(2 downto 0);                     -- awprot
			h2f_lw_AWVALID           : out   std_logic;                                        -- awvalid
			h2f_lw_AWREADY           : in    std_logic                     := 'X';             -- awready
			h2f_lw_WID               : out   std_logic_vector(11 downto 0);                    -- wid
			h2f_lw_WDATA             : out   std_logic_vector(31 downto 0);                    -- wdata
			h2f_lw_WSTRB             : out   std_logic_vector(3 downto 0);                     -- wstrb
			h2f_lw_WLAST             : out   std_logic;                                        -- wlast
			h2f_lw_WVALID            : out   std_logic;                                        -- wvalid
			h2f_lw_WREADY            : in    std_logic                     := 'X';             -- wready
			h2f_lw_BID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- bid
			h2f_lw_BRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- bresp
			h2f_lw_BVALID            : in    std_logic                     := 'X';             -- bvalid
			h2f_lw_BREADY            : out   std_logic;                                        -- bready
			h2f_lw_ARID              : out   std_logic_vector(11 downto 0);                    -- arid
			h2f_lw_ARADDR            : out   std_logic_vector(20 downto 0);                    -- araddr
			h2f_lw_ARLEN             : out   std_logic_vector(3 downto 0);                     -- arlen
			h2f_lw_ARSIZE            : out   std_logic_vector(2 downto 0);                     -- arsize
			h2f_lw_ARBURST           : out   std_logic_vector(1 downto 0);                     -- arburst
			h2f_lw_ARLOCK            : out   std_logic_vector(1 downto 0);                     -- arlock
			h2f_lw_ARCACHE           : out   std_logic_vector(3 downto 0);                     -- arcache
			h2f_lw_ARPROT            : out   std_logic_vector(2 downto 0);                     -- arprot
			h2f_lw_ARVALID           : out   std_logic;                                        -- arvalid
			h2f_lw_ARREADY           : in    std_logic                     := 'X';             -- arready
			h2f_lw_RID               : in    std_logic_vector(11 downto 0) := (others => 'X'); -- rid
			h2f_lw_RDATA             : in    std_logic_vector(31 downto 0) := (others => 'X'); -- rdata
			h2f_lw_RRESP             : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- rresp
			h2f_lw_RLAST             : in    std_logic                     := 'X';             -- rlast
			h2f_lw_RVALID            : in    std_logic                     := 'X';             -- rvalid
			h2f_lw_RREADY            : out   std_logic                                         -- rready
		);
	end component soc_system_hps_0;

	component soc_system_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component soc_system_sysid_qsys_0;

	component soc_system_mm_interconnect_0 is
		port (
			hps_0_h2f_lw_axi_master_awid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- awid
			hps_0_h2f_lw_axi_master_awaddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- awaddr
			hps_0_h2f_lw_axi_master_awlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awlen
			hps_0_h2f_lw_axi_master_awsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awsize
			hps_0_h2f_lw_axi_master_awburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awburst
			hps_0_h2f_lw_axi_master_awlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- awlock
			hps_0_h2f_lw_axi_master_awcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- awcache
			hps_0_h2f_lw_axi_master_awprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- awprot
			hps_0_h2f_lw_axi_master_awvalid                                     : in  std_logic                     := 'X';             -- awvalid
			hps_0_h2f_lw_axi_master_awready                                     : out std_logic;                                        -- awready
			hps_0_h2f_lw_axi_master_wid                                         : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wid
			hps_0_h2f_lw_axi_master_wdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wdata
			hps_0_h2f_lw_axi_master_wstrb                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wstrb
			hps_0_h2f_lw_axi_master_wlast                                       : in  std_logic                     := 'X';             -- wlast
			hps_0_h2f_lw_axi_master_wvalid                                      : in  std_logic                     := 'X';             -- wvalid
			hps_0_h2f_lw_axi_master_wready                                      : out std_logic;                                        -- wready
			hps_0_h2f_lw_axi_master_bid                                         : out std_logic_vector(11 downto 0);                    -- bid
			hps_0_h2f_lw_axi_master_bresp                                       : out std_logic_vector(1 downto 0);                     -- bresp
			hps_0_h2f_lw_axi_master_bvalid                                      : out std_logic;                                        -- bvalid
			hps_0_h2f_lw_axi_master_bready                                      : in  std_logic                     := 'X';             -- bready
			hps_0_h2f_lw_axi_master_arid                                        : in  std_logic_vector(11 downto 0) := (others => 'X'); -- arid
			hps_0_h2f_lw_axi_master_araddr                                      : in  std_logic_vector(20 downto 0) := (others => 'X'); -- araddr
			hps_0_h2f_lw_axi_master_arlen                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arlen
			hps_0_h2f_lw_axi_master_arsize                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arsize
			hps_0_h2f_lw_axi_master_arburst                                     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arburst
			hps_0_h2f_lw_axi_master_arlock                                      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- arlock
			hps_0_h2f_lw_axi_master_arcache                                     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- arcache
			hps_0_h2f_lw_axi_master_arprot                                      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- arprot
			hps_0_h2f_lw_axi_master_arvalid                                     : in  std_logic                     := 'X';             -- arvalid
			hps_0_h2f_lw_axi_master_arready                                     : out std_logic;                                        -- arready
			hps_0_h2f_lw_axi_master_rid                                         : out std_logic_vector(11 downto 0);                    -- rid
			hps_0_h2f_lw_axi_master_rdata                                       : out std_logic_vector(31 downto 0);                    -- rdata
			hps_0_h2f_lw_axi_master_rresp                                       : out std_logic_vector(1 downto 0);                     -- rresp
			hps_0_h2f_lw_axi_master_rlast                                       : out std_logic;                                        -- rlast
			hps_0_h2f_lw_axi_master_rvalid                                      : out std_logic;                                        -- rvalid
			hps_0_h2f_lw_axi_master_rready                                      : in  std_logic                     := 'X';             -- rready
			clk_0_clk_clk                                                       : in  std_logic                     := 'X';             -- clk
			Easy_Driver_Y_reset_reset_bridge_in_reset_reset                     : in  std_logic                     := 'X';             -- reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			Easy_Driver_X_avalon_slave_dir_write                                : out std_logic;                                        -- write
			Easy_Driver_X_avalon_slave_dir_read                                 : out std_logic;                                        -- read
			Easy_Driver_X_avalon_slave_dir_readdata                             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			Easy_Driver_X_avalon_slave_dir_writedata                            : out std_logic_vector(7 downto 0);                     -- writedata
			Easy_Driver_X_avalon_slave_duty_write                               : out std_logic;                                        -- write
			Easy_Driver_X_avalon_slave_duty_read                                : out std_logic;                                        -- read
			Easy_Driver_X_avalon_slave_duty_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Easy_Driver_X_avalon_slave_duty_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			Easy_Driver_X_avalon_slave_period_write                             : out std_logic;                                        -- write
			Easy_Driver_X_avalon_slave_period_read                              : out std_logic;                                        -- read
			Easy_Driver_X_avalon_slave_period_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Easy_Driver_X_avalon_slave_period_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			Easy_Driver_X_avalon_slave_step_write                               : out std_logic;                                        -- write
			Easy_Driver_X_avalon_slave_step_read                                : out std_logic;                                        -- read
			Easy_Driver_X_avalon_slave_step_readdata                            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Easy_Driver_X_avalon_slave_step_writedata                           : out std_logic_vector(15 downto 0);                    -- writedata
			Easy_Driver_Y_avalon_slave_dir_write                                : out std_logic;                                        -- write
			Easy_Driver_Y_avalon_slave_dir_read                                 : out std_logic;                                        -- read
			Easy_Driver_Y_avalon_slave_dir_readdata                             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			Easy_Driver_Y_avalon_slave_dir_writedata                            : out std_logic_vector(7 downto 0);                     -- writedata
			Easy_Driver_Y_avalon_slave_duty_write                               : out std_logic;                                        -- write
			Easy_Driver_Y_avalon_slave_duty_read                                : out std_logic;                                        -- read
			Easy_Driver_Y_avalon_slave_duty_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Easy_Driver_Y_avalon_slave_duty_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			Easy_Driver_Y_avalon_slave_period_write                             : out std_logic;                                        -- write
			Easy_Driver_Y_avalon_slave_period_read                              : out std_logic;                                        -- read
			Easy_Driver_Y_avalon_slave_period_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			Easy_Driver_Y_avalon_slave_period_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			Easy_Driver_Y_avalon_slave_step_write                               : out std_logic;                                        -- write
			Easy_Driver_Y_avalon_slave_step_read                                : out std_logic;                                        -- read
			Easy_Driver_Y_avalon_slave_step_readdata                            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			Easy_Driver_Y_avalon_slave_step_writedata                           : out std_logic_vector(15 downto 0);                    -- writedata
			sysid_qsys_0_control_slave_address                                  : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component soc_system_mm_interconnect_0;

	component soc_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller;

	component soc_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component soc_system_rst_controller_001;

	signal hps_0_h2f_lw_axi_master_awburst                                     : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	signal hps_0_h2f_lw_axi_master_arlen                                       : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	signal hps_0_h2f_lw_axi_master_wstrb                                       : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	signal hps_0_h2f_lw_axi_master_wready                                      : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	signal hps_0_h2f_lw_axi_master_rid                                         : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	signal hps_0_h2f_lw_axi_master_rready                                      : std_logic;                     -- hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	signal hps_0_h2f_lw_axi_master_awlen                                       : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	signal hps_0_h2f_lw_axi_master_wid                                         : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	signal hps_0_h2f_lw_axi_master_arcache                                     : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	signal hps_0_h2f_lw_axi_master_wvalid                                      : std_logic;                     -- hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	signal hps_0_h2f_lw_axi_master_araddr                                      : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	signal hps_0_h2f_lw_axi_master_arprot                                      : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	signal hps_0_h2f_lw_axi_master_awprot                                      : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	signal hps_0_h2f_lw_axi_master_wdata                                       : std_logic_vector(31 downto 0); -- hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	signal hps_0_h2f_lw_axi_master_arvalid                                     : std_logic;                     -- hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	signal hps_0_h2f_lw_axi_master_awcache                                     : std_logic_vector(3 downto 0);  -- hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	signal hps_0_h2f_lw_axi_master_arid                                        : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	signal hps_0_h2f_lw_axi_master_arlock                                      : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	signal hps_0_h2f_lw_axi_master_awlock                                      : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	signal hps_0_h2f_lw_axi_master_awaddr                                      : std_logic_vector(20 downto 0); -- hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	signal hps_0_h2f_lw_axi_master_bresp                                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	signal hps_0_h2f_lw_axi_master_arready                                     : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	signal hps_0_h2f_lw_axi_master_rdata                                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	signal hps_0_h2f_lw_axi_master_awready                                     : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	signal hps_0_h2f_lw_axi_master_arburst                                     : std_logic_vector(1 downto 0);  -- hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	signal hps_0_h2f_lw_axi_master_arsize                                      : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	signal hps_0_h2f_lw_axi_master_bready                                      : std_logic;                     -- hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	signal hps_0_h2f_lw_axi_master_rlast                                       : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	signal hps_0_h2f_lw_axi_master_wlast                                       : std_logic;                     -- hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	signal hps_0_h2f_lw_axi_master_rresp                                       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	signal hps_0_h2f_lw_axi_master_awid                                        : std_logic_vector(11 downto 0); -- hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	signal hps_0_h2f_lw_axi_master_bid                                         : std_logic_vector(11 downto 0); -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	signal hps_0_h2f_lw_axi_master_bvalid                                      : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	signal hps_0_h2f_lw_axi_master_awsize                                      : std_logic_vector(2 downto 0);  -- hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	signal hps_0_h2f_lw_axi_master_awvalid                                     : std_logic;                     -- hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	signal hps_0_h2f_lw_axi_master_rvalid                                      : std_logic;                     -- mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	signal mm_interconnect_0_easy_driver_y_avalon_slave_dir_readdata           : std_logic_vector(7 downto 0);  -- Easy_Driver_Y:dir_readdata -> mm_interconnect_0:Easy_Driver_Y_avalon_slave_dir_readdata
	signal mm_interconnect_0_easy_driver_y_avalon_slave_dir_read               : std_logic;                     -- mm_interconnect_0:Easy_Driver_Y_avalon_slave_dir_read -> mm_interconnect_0_easy_driver_y_avalon_slave_dir_read:in
	signal mm_interconnect_0_easy_driver_y_avalon_slave_dir_write              : std_logic;                     -- mm_interconnect_0:Easy_Driver_Y_avalon_slave_dir_write -> mm_interconnect_0_easy_driver_y_avalon_slave_dir_write:in
	signal mm_interconnect_0_easy_driver_y_avalon_slave_dir_writedata          : std_logic_vector(7 downto 0);  -- mm_interconnect_0:Easy_Driver_Y_avalon_slave_dir_writedata -> Easy_Driver_Y:dir_writedata
	signal mm_interconnect_0_easy_driver_x_avalon_slave_dir_readdata           : std_logic_vector(7 downto 0);  -- Easy_Driver_X:dir_readdata -> mm_interconnect_0:Easy_Driver_X_avalon_slave_dir_readdata
	signal mm_interconnect_0_easy_driver_x_avalon_slave_dir_read               : std_logic;                     -- mm_interconnect_0:Easy_Driver_X_avalon_slave_dir_read -> mm_interconnect_0_easy_driver_x_avalon_slave_dir_read:in
	signal mm_interconnect_0_easy_driver_x_avalon_slave_dir_write              : std_logic;                     -- mm_interconnect_0:Easy_Driver_X_avalon_slave_dir_write -> mm_interconnect_0_easy_driver_x_avalon_slave_dir_write:in
	signal mm_interconnect_0_easy_driver_x_avalon_slave_dir_writedata          : std_logic_vector(7 downto 0);  -- mm_interconnect_0:Easy_Driver_X_avalon_slave_dir_writedata -> Easy_Driver_X:dir_writedata
	signal mm_interconnect_0_easy_driver_y_avalon_slave_duty_readdata          : std_logic_vector(31 downto 0); -- Easy_Driver_Y:duty_readdata -> mm_interconnect_0:Easy_Driver_Y_avalon_slave_duty_readdata
	signal mm_interconnect_0_easy_driver_y_avalon_slave_duty_read              : std_logic;                     -- mm_interconnect_0:Easy_Driver_Y_avalon_slave_duty_read -> mm_interconnect_0_easy_driver_y_avalon_slave_duty_read:in
	signal mm_interconnect_0_easy_driver_y_avalon_slave_duty_write             : std_logic;                     -- mm_interconnect_0:Easy_Driver_Y_avalon_slave_duty_write -> mm_interconnect_0_easy_driver_y_avalon_slave_duty_write:in
	signal mm_interconnect_0_easy_driver_y_avalon_slave_duty_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:Easy_Driver_Y_avalon_slave_duty_writedata -> Easy_Driver_Y:duty_writedata
	signal mm_interconnect_0_easy_driver_x_avalon_slave_duty_readdata          : std_logic_vector(31 downto 0); -- Easy_Driver_X:duty_readdata -> mm_interconnect_0:Easy_Driver_X_avalon_slave_duty_readdata
	signal mm_interconnect_0_easy_driver_x_avalon_slave_duty_read              : std_logic;                     -- mm_interconnect_0:Easy_Driver_X_avalon_slave_duty_read -> mm_interconnect_0_easy_driver_x_avalon_slave_duty_read:in
	signal mm_interconnect_0_easy_driver_x_avalon_slave_duty_write             : std_logic;                     -- mm_interconnect_0:Easy_Driver_X_avalon_slave_duty_write -> mm_interconnect_0_easy_driver_x_avalon_slave_duty_write:in
	signal mm_interconnect_0_easy_driver_x_avalon_slave_duty_writedata         : std_logic_vector(31 downto 0); -- mm_interconnect_0:Easy_Driver_X_avalon_slave_duty_writedata -> Easy_Driver_X:duty_writedata
	signal mm_interconnect_0_easy_driver_y_avalon_slave_period_readdata        : std_logic_vector(31 downto 0); -- Easy_Driver_Y:period_readdata -> mm_interconnect_0:Easy_Driver_Y_avalon_slave_period_readdata
	signal mm_interconnect_0_easy_driver_y_avalon_slave_period_read            : std_logic;                     -- mm_interconnect_0:Easy_Driver_Y_avalon_slave_period_read -> mm_interconnect_0_easy_driver_y_avalon_slave_period_read:in
	signal mm_interconnect_0_easy_driver_y_avalon_slave_period_write           : std_logic;                     -- mm_interconnect_0:Easy_Driver_Y_avalon_slave_period_write -> mm_interconnect_0_easy_driver_y_avalon_slave_period_write:in
	signal mm_interconnect_0_easy_driver_y_avalon_slave_period_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:Easy_Driver_Y_avalon_slave_period_writedata -> Easy_Driver_Y:period_writedata
	signal mm_interconnect_0_easy_driver_x_avalon_slave_period_readdata        : std_logic_vector(31 downto 0); -- Easy_Driver_X:period_readdata -> mm_interconnect_0:Easy_Driver_X_avalon_slave_period_readdata
	signal mm_interconnect_0_easy_driver_x_avalon_slave_period_read            : std_logic;                     -- mm_interconnect_0:Easy_Driver_X_avalon_slave_period_read -> mm_interconnect_0_easy_driver_x_avalon_slave_period_read:in
	signal mm_interconnect_0_easy_driver_x_avalon_slave_period_write           : std_logic;                     -- mm_interconnect_0:Easy_Driver_X_avalon_slave_period_write -> mm_interconnect_0_easy_driver_x_avalon_slave_period_write:in
	signal mm_interconnect_0_easy_driver_x_avalon_slave_period_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:Easy_Driver_X_avalon_slave_period_writedata -> Easy_Driver_X:period_writedata
	signal mm_interconnect_0_easy_driver_y_avalon_slave_step_readdata          : std_logic_vector(15 downto 0); -- Easy_Driver_Y:step_readdata -> mm_interconnect_0:Easy_Driver_Y_avalon_slave_step_readdata
	signal mm_interconnect_0_easy_driver_y_avalon_slave_step_read              : std_logic;                     -- mm_interconnect_0:Easy_Driver_Y_avalon_slave_step_read -> mm_interconnect_0_easy_driver_y_avalon_slave_step_read:in
	signal mm_interconnect_0_easy_driver_y_avalon_slave_step_write             : std_logic;                     -- mm_interconnect_0:Easy_Driver_Y_avalon_slave_step_write -> mm_interconnect_0_easy_driver_y_avalon_slave_step_write:in
	signal mm_interconnect_0_easy_driver_y_avalon_slave_step_writedata         : std_logic_vector(15 downto 0); -- mm_interconnect_0:Easy_Driver_Y_avalon_slave_step_writedata -> Easy_Driver_Y:step_writedata
	signal mm_interconnect_0_easy_driver_x_avalon_slave_step_readdata          : std_logic_vector(15 downto 0); -- Easy_Driver_X:step_readdata -> mm_interconnect_0:Easy_Driver_X_avalon_slave_step_readdata
	signal mm_interconnect_0_easy_driver_x_avalon_slave_step_read              : std_logic;                     -- mm_interconnect_0:Easy_Driver_X_avalon_slave_step_read -> mm_interconnect_0_easy_driver_x_avalon_slave_step_read:in
	signal mm_interconnect_0_easy_driver_x_avalon_slave_step_write             : std_logic;                     -- mm_interconnect_0:Easy_Driver_X_avalon_slave_step_write -> mm_interconnect_0_easy_driver_x_avalon_slave_step_write:in
	signal mm_interconnect_0_easy_driver_x_avalon_slave_step_writedata         : std_logic_vector(15 downto 0); -- mm_interconnect_0:Easy_Driver_X_avalon_slave_step_writedata -> Easy_Driver_X:step_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata               : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address                : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal rst_controller_reset_out_reset                                      : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:Easy_Driver_Y_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal hps_0_h2f_reset_reset                                               : std_logic;                     -- hps_0:h2f_rst_n -> hps_0_h2f_reset_reset:in
	signal rst_controller_001_reset_out_reset                                  : std_logic;                     -- rst_controller_001:reset_out -> mm_interconnect_0:hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset
	signal reset_reset_n_ports_inv                                             : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_easy_driver_y_avalon_slave_dir_read_ports_inv     : std_logic;                     -- mm_interconnect_0_easy_driver_y_avalon_slave_dir_read:inv -> Easy_Driver_Y:dir_read_n
	signal mm_interconnect_0_easy_driver_y_avalon_slave_dir_write_ports_inv    : std_logic;                     -- mm_interconnect_0_easy_driver_y_avalon_slave_dir_write:inv -> Easy_Driver_Y:dir_write_n
	signal mm_interconnect_0_easy_driver_x_avalon_slave_dir_read_ports_inv     : std_logic;                     -- mm_interconnect_0_easy_driver_x_avalon_slave_dir_read:inv -> Easy_Driver_X:dir_read_n
	signal mm_interconnect_0_easy_driver_x_avalon_slave_dir_write_ports_inv    : std_logic;                     -- mm_interconnect_0_easy_driver_x_avalon_slave_dir_write:inv -> Easy_Driver_X:dir_write_n
	signal mm_interconnect_0_easy_driver_y_avalon_slave_duty_read_ports_inv    : std_logic;                     -- mm_interconnect_0_easy_driver_y_avalon_slave_duty_read:inv -> Easy_Driver_Y:duty_read_n
	signal mm_interconnect_0_easy_driver_y_avalon_slave_duty_write_ports_inv   : std_logic;                     -- mm_interconnect_0_easy_driver_y_avalon_slave_duty_write:inv -> Easy_Driver_Y:duty_write_n
	signal mm_interconnect_0_easy_driver_x_avalon_slave_duty_read_ports_inv    : std_logic;                     -- mm_interconnect_0_easy_driver_x_avalon_slave_duty_read:inv -> Easy_Driver_X:duty_read_n
	signal mm_interconnect_0_easy_driver_x_avalon_slave_duty_write_ports_inv   : std_logic;                     -- mm_interconnect_0_easy_driver_x_avalon_slave_duty_write:inv -> Easy_Driver_X:duty_write_n
	signal mm_interconnect_0_easy_driver_y_avalon_slave_period_read_ports_inv  : std_logic;                     -- mm_interconnect_0_easy_driver_y_avalon_slave_period_read:inv -> Easy_Driver_Y:period_read_n
	signal mm_interconnect_0_easy_driver_y_avalon_slave_period_write_ports_inv : std_logic;                     -- mm_interconnect_0_easy_driver_y_avalon_slave_period_write:inv -> Easy_Driver_Y:period_write_n
	signal mm_interconnect_0_easy_driver_x_avalon_slave_period_read_ports_inv  : std_logic;                     -- mm_interconnect_0_easy_driver_x_avalon_slave_period_read:inv -> Easy_Driver_X:period_read_n
	signal mm_interconnect_0_easy_driver_x_avalon_slave_period_write_ports_inv : std_logic;                     -- mm_interconnect_0_easy_driver_x_avalon_slave_period_write:inv -> Easy_Driver_X:period_write_n
	signal mm_interconnect_0_easy_driver_y_avalon_slave_step_read_ports_inv    : std_logic;                     -- mm_interconnect_0_easy_driver_y_avalon_slave_step_read:inv -> Easy_Driver_Y:step_read_n
	signal mm_interconnect_0_easy_driver_y_avalon_slave_step_write_ports_inv   : std_logic;                     -- mm_interconnect_0_easy_driver_y_avalon_slave_step_write:inv -> Easy_Driver_Y:step_write_n
	signal mm_interconnect_0_easy_driver_x_avalon_slave_step_read_ports_inv    : std_logic;                     -- mm_interconnect_0_easy_driver_x_avalon_slave_step_read:inv -> Easy_Driver_X:step_read_n
	signal mm_interconnect_0_easy_driver_x_avalon_slave_step_write_ports_inv   : std_logic;                     -- mm_interconnect_0_easy_driver_x_avalon_slave_step_write:inv -> Easy_Driver_X:step_write_n
	signal rst_controller_reset_out_reset_ports_inv                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [Easy_Driver_X:reset_n, Easy_Driver_Y:reset_n, sysid_qsys_0:reset_n]
	signal hps_0_h2f_reset_reset_ports_inv                                     : std_logic;                     -- hps_0_h2f_reset_reset:inv -> [rst_controller:reset_in1, rst_controller_001:reset_in0]

begin

	easy_driver_x : component Easy_Driver
		port map (
			clk                => clk_clk,                                                             --               clock.clk
			reset_n            => rst_controller_reset_out_reset_ports_inv,                            --               reset.reset_n
			conduit_end_dir    => easy_driver_x_conduit_end_dir,                                       --         conduit_end.dir
			conduit_end_step   => easy_driver_x_conduit_end_step,                                      --                    .step
			conduit_end_enable => easy_driver_x_conduit_end_enable,                                    --                    .enable
			step_read_n        => mm_interconnect_0_easy_driver_x_avalon_slave_step_read_ports_inv,    --   avalon_slave_step.read_n
			step_readdata      => mm_interconnect_0_easy_driver_x_avalon_slave_step_readdata,          --                    .readdata
			step_write_n       => mm_interconnect_0_easy_driver_x_avalon_slave_step_write_ports_inv,   --                    .write_n
			step_writedata     => mm_interconnect_0_easy_driver_x_avalon_slave_step_writedata,         --                    .writedata
			dir_read_n         => mm_interconnect_0_easy_driver_x_avalon_slave_dir_read_ports_inv,     --    avalon_slave_dir.read_n
			dir_readdata       => mm_interconnect_0_easy_driver_x_avalon_slave_dir_readdata,           --                    .readdata
			dir_write_n        => mm_interconnect_0_easy_driver_x_avalon_slave_dir_write_ports_inv,    --                    .write_n
			dir_writedata      => mm_interconnect_0_easy_driver_x_avalon_slave_dir_writedata,          --                    .writedata
			period_read_n      => mm_interconnect_0_easy_driver_x_avalon_slave_period_read_ports_inv,  -- avalon_slave_period.read_n
			period_readdata    => mm_interconnect_0_easy_driver_x_avalon_slave_period_readdata,        --                    .readdata
			period_write_n     => mm_interconnect_0_easy_driver_x_avalon_slave_period_write_ports_inv, --                    .write_n
			period_writedata   => mm_interconnect_0_easy_driver_x_avalon_slave_period_writedata,       --                    .writedata
			duty_read_n        => mm_interconnect_0_easy_driver_x_avalon_slave_duty_read_ports_inv,    --   avalon_slave_duty.read_n
			duty_readdata      => mm_interconnect_0_easy_driver_x_avalon_slave_duty_readdata,          --                    .readdata
			duty_write_n       => mm_interconnect_0_easy_driver_x_avalon_slave_duty_write_ports_inv,   --                    .write_n
			duty_writedata     => mm_interconnect_0_easy_driver_x_avalon_slave_duty_writedata          --                    .writedata
		);

	easy_driver_y : component Easy_Driver
		port map (
			clk                => clk_clk,                                                             --               clock.clk
			reset_n            => rst_controller_reset_out_reset_ports_inv,                            --               reset.reset_n
			conduit_end_dir    => easy_driver_y_conduit_end_dir,                                       --         conduit_end.dir
			conduit_end_step   => easy_driver_y_conduit_end_step,                                      --                    .step
			conduit_end_enable => easy_driver_y_conduit_end_enable,                                    --                    .enable
			step_read_n        => mm_interconnect_0_easy_driver_y_avalon_slave_step_read_ports_inv,    --   avalon_slave_step.read_n
			step_readdata      => mm_interconnect_0_easy_driver_y_avalon_slave_step_readdata,          --                    .readdata
			step_write_n       => mm_interconnect_0_easy_driver_y_avalon_slave_step_write_ports_inv,   --                    .write_n
			step_writedata     => mm_interconnect_0_easy_driver_y_avalon_slave_step_writedata,         --                    .writedata
			dir_read_n         => mm_interconnect_0_easy_driver_y_avalon_slave_dir_read_ports_inv,     --    avalon_slave_dir.read_n
			dir_readdata       => mm_interconnect_0_easy_driver_y_avalon_slave_dir_readdata,           --                    .readdata
			dir_write_n        => mm_interconnect_0_easy_driver_y_avalon_slave_dir_write_ports_inv,    --                    .write_n
			dir_writedata      => mm_interconnect_0_easy_driver_y_avalon_slave_dir_writedata,          --                    .writedata
			period_read_n      => mm_interconnect_0_easy_driver_y_avalon_slave_period_read_ports_inv,  -- avalon_slave_period.read_n
			period_readdata    => mm_interconnect_0_easy_driver_y_avalon_slave_period_readdata,        --                    .readdata
			period_write_n     => mm_interconnect_0_easy_driver_y_avalon_slave_period_write_ports_inv, --                    .write_n
			period_writedata   => mm_interconnect_0_easy_driver_y_avalon_slave_period_writedata,       --                    .writedata
			duty_read_n        => mm_interconnect_0_easy_driver_y_avalon_slave_duty_read_ports_inv,    --   avalon_slave_duty.read_n
			duty_readdata      => mm_interconnect_0_easy_driver_y_avalon_slave_duty_readdata,          --                    .readdata
			duty_write_n       => mm_interconnect_0_easy_driver_y_avalon_slave_duty_write_ports_inv,   --                    .write_n
			duty_writedata     => mm_interconnect_0_easy_driver_y_avalon_slave_duty_writedata          --                    .writedata
		);

	hps_0 : component soc_system_hps_0
		generic map (
			F2S_Width => 0,
			S2F_Width => 0
		)
		port map (
			mem_a                    => memory_mem_a,                    --            memory.mem_a
			mem_ba                   => memory_mem_ba,                   --                  .mem_ba
			mem_ck                   => memory_mem_ck,                   --                  .mem_ck
			mem_ck_n                 => memory_mem_ck_n,                 --                  .mem_ck_n
			mem_cke                  => memory_mem_cke,                  --                  .mem_cke
			mem_cs_n                 => memory_mem_cs_n,                 --                  .mem_cs_n
			mem_ras_n                => memory_mem_ras_n,                --                  .mem_ras_n
			mem_cas_n                => memory_mem_cas_n,                --                  .mem_cas_n
			mem_we_n                 => memory_mem_we_n,                 --                  .mem_we_n
			mem_reset_n              => memory_mem_reset_n,              --                  .mem_reset_n
			mem_dq                   => memory_mem_dq,                   --                  .mem_dq
			mem_dqs                  => memory_mem_dqs,                  --                  .mem_dqs
			mem_dqs_n                => memory_mem_dqs_n,                --                  .mem_dqs_n
			mem_odt                  => memory_mem_odt,                  --                  .mem_odt
			mem_dm                   => memory_mem_dm,                   --                  .mem_dm
			oct_rzqin                => memory_oct_rzqin,                --                  .oct_rzqin
			hps_io_emac1_inst_TX_CLK => hps_io_hps_io_emac1_inst_TX_CLK, --            hps_io.hps_io_emac1_inst_TX_CLK
			hps_io_emac1_inst_TXD0   => hps_io_hps_io_emac1_inst_TXD0,   --                  .hps_io_emac1_inst_TXD0
			hps_io_emac1_inst_TXD1   => hps_io_hps_io_emac1_inst_TXD1,   --                  .hps_io_emac1_inst_TXD1
			hps_io_emac1_inst_TXD2   => hps_io_hps_io_emac1_inst_TXD2,   --                  .hps_io_emac1_inst_TXD2
			hps_io_emac1_inst_TXD3   => hps_io_hps_io_emac1_inst_TXD3,   --                  .hps_io_emac1_inst_TXD3
			hps_io_emac1_inst_RXD0   => hps_io_hps_io_emac1_inst_RXD0,   --                  .hps_io_emac1_inst_RXD0
			hps_io_emac1_inst_MDIO   => hps_io_hps_io_emac1_inst_MDIO,   --                  .hps_io_emac1_inst_MDIO
			hps_io_emac1_inst_MDC    => hps_io_hps_io_emac1_inst_MDC,    --                  .hps_io_emac1_inst_MDC
			hps_io_emac1_inst_RX_CTL => hps_io_hps_io_emac1_inst_RX_CTL, --                  .hps_io_emac1_inst_RX_CTL
			hps_io_emac1_inst_TX_CTL => hps_io_hps_io_emac1_inst_TX_CTL, --                  .hps_io_emac1_inst_TX_CTL
			hps_io_emac1_inst_RX_CLK => hps_io_hps_io_emac1_inst_RX_CLK, --                  .hps_io_emac1_inst_RX_CLK
			hps_io_emac1_inst_RXD1   => hps_io_hps_io_emac1_inst_RXD1,   --                  .hps_io_emac1_inst_RXD1
			hps_io_emac1_inst_RXD2   => hps_io_hps_io_emac1_inst_RXD2,   --                  .hps_io_emac1_inst_RXD2
			hps_io_emac1_inst_RXD3   => hps_io_hps_io_emac1_inst_RXD3,   --                  .hps_io_emac1_inst_RXD3
			hps_io_sdio_inst_CMD     => hps_io_hps_io_sdio_inst_CMD,     --                  .hps_io_sdio_inst_CMD
			hps_io_sdio_inst_D0      => hps_io_hps_io_sdio_inst_D0,      --                  .hps_io_sdio_inst_D0
			hps_io_sdio_inst_D1      => hps_io_hps_io_sdio_inst_D1,      --                  .hps_io_sdio_inst_D1
			hps_io_sdio_inst_CLK     => hps_io_hps_io_sdio_inst_CLK,     --                  .hps_io_sdio_inst_CLK
			hps_io_sdio_inst_D2      => hps_io_hps_io_sdio_inst_D2,      --                  .hps_io_sdio_inst_D2
			hps_io_sdio_inst_D3      => hps_io_hps_io_sdio_inst_D3,      --                  .hps_io_sdio_inst_D3
			hps_io_usb1_inst_D0      => hps_io_hps_io_usb1_inst_D0,      --                  .hps_io_usb1_inst_D0
			hps_io_usb1_inst_D1      => hps_io_hps_io_usb1_inst_D1,      --                  .hps_io_usb1_inst_D1
			hps_io_usb1_inst_D2      => hps_io_hps_io_usb1_inst_D2,      --                  .hps_io_usb1_inst_D2
			hps_io_usb1_inst_D3      => hps_io_hps_io_usb1_inst_D3,      --                  .hps_io_usb1_inst_D3
			hps_io_usb1_inst_D4      => hps_io_hps_io_usb1_inst_D4,      --                  .hps_io_usb1_inst_D4
			hps_io_usb1_inst_D5      => hps_io_hps_io_usb1_inst_D5,      --                  .hps_io_usb1_inst_D5
			hps_io_usb1_inst_D6      => hps_io_hps_io_usb1_inst_D6,      --                  .hps_io_usb1_inst_D6
			hps_io_usb1_inst_D7      => hps_io_hps_io_usb1_inst_D7,      --                  .hps_io_usb1_inst_D7
			hps_io_usb1_inst_CLK     => hps_io_hps_io_usb1_inst_CLK,     --                  .hps_io_usb1_inst_CLK
			hps_io_usb1_inst_STP     => hps_io_hps_io_usb1_inst_STP,     --                  .hps_io_usb1_inst_STP
			hps_io_usb1_inst_DIR     => hps_io_hps_io_usb1_inst_DIR,     --                  .hps_io_usb1_inst_DIR
			hps_io_usb1_inst_NXT     => hps_io_hps_io_usb1_inst_NXT,     --                  .hps_io_usb1_inst_NXT
			hps_io_spim1_inst_CLK    => hps_io_hps_io_spim1_inst_CLK,    --                  .hps_io_spim1_inst_CLK
			hps_io_spim1_inst_MOSI   => hps_io_hps_io_spim1_inst_MOSI,   --                  .hps_io_spim1_inst_MOSI
			hps_io_spim1_inst_MISO   => hps_io_hps_io_spim1_inst_MISO,   --                  .hps_io_spim1_inst_MISO
			hps_io_spim1_inst_SS0    => hps_io_hps_io_spim1_inst_SS0,    --                  .hps_io_spim1_inst_SS0
			hps_io_uart0_inst_RX     => hps_io_hps_io_uart0_inst_RX,     --                  .hps_io_uart0_inst_RX
			hps_io_uart0_inst_TX     => hps_io_hps_io_uart0_inst_TX,     --                  .hps_io_uart0_inst_TX
			hps_io_i2c0_inst_SDA     => hps_io_hps_io_i2c0_inst_SDA,     --                  .hps_io_i2c0_inst_SDA
			hps_io_i2c0_inst_SCL     => hps_io_hps_io_i2c0_inst_SCL,     --                  .hps_io_i2c0_inst_SCL
			hps_io_i2c1_inst_SDA     => hps_io_hps_io_i2c1_inst_SDA,     --                  .hps_io_i2c1_inst_SDA
			hps_io_i2c1_inst_SCL     => hps_io_hps_io_i2c1_inst_SCL,     --                  .hps_io_i2c1_inst_SCL
			hps_io_gpio_inst_GPIO09  => hps_io_hps_io_gpio_inst_GPIO09,  --                  .hps_io_gpio_inst_GPIO09
			hps_io_gpio_inst_GPIO35  => hps_io_hps_io_gpio_inst_GPIO35,  --                  .hps_io_gpio_inst_GPIO35
			hps_io_gpio_inst_GPIO40  => hps_io_hps_io_gpio_inst_GPIO40,  --                  .hps_io_gpio_inst_GPIO40
			hps_io_gpio_inst_GPIO48  => hps_io_hps_io_gpio_inst_GPIO48,  --                  .hps_io_gpio_inst_GPIO48
			hps_io_gpio_inst_GPIO53  => hps_io_hps_io_gpio_inst_GPIO53,  --                  .hps_io_gpio_inst_GPIO53
			hps_io_gpio_inst_GPIO54  => hps_io_hps_io_gpio_inst_GPIO54,  --                  .hps_io_gpio_inst_GPIO54
			hps_io_gpio_inst_GPIO61  => hps_io_hps_io_gpio_inst_GPIO61,  --                  .hps_io_gpio_inst_GPIO61
			h2f_rst_n                => hps_0_h2f_reset_reset,           --         h2f_reset.reset_n
			h2f_lw_axi_clk           => clk_clk,                         --  h2f_lw_axi_clock.clk
			h2f_lw_AWID              => hps_0_h2f_lw_axi_master_awid,    -- h2f_lw_axi_master.awid
			h2f_lw_AWADDR            => hps_0_h2f_lw_axi_master_awaddr,  --                  .awaddr
			h2f_lw_AWLEN             => hps_0_h2f_lw_axi_master_awlen,   --                  .awlen
			h2f_lw_AWSIZE            => hps_0_h2f_lw_axi_master_awsize,  --                  .awsize
			h2f_lw_AWBURST           => hps_0_h2f_lw_axi_master_awburst, --                  .awburst
			h2f_lw_AWLOCK            => hps_0_h2f_lw_axi_master_awlock,  --                  .awlock
			h2f_lw_AWCACHE           => hps_0_h2f_lw_axi_master_awcache, --                  .awcache
			h2f_lw_AWPROT            => hps_0_h2f_lw_axi_master_awprot,  --                  .awprot
			h2f_lw_AWVALID           => hps_0_h2f_lw_axi_master_awvalid, --                  .awvalid
			h2f_lw_AWREADY           => hps_0_h2f_lw_axi_master_awready, --                  .awready
			h2f_lw_WID               => hps_0_h2f_lw_axi_master_wid,     --                  .wid
			h2f_lw_WDATA             => hps_0_h2f_lw_axi_master_wdata,   --                  .wdata
			h2f_lw_WSTRB             => hps_0_h2f_lw_axi_master_wstrb,   --                  .wstrb
			h2f_lw_WLAST             => hps_0_h2f_lw_axi_master_wlast,   --                  .wlast
			h2f_lw_WVALID            => hps_0_h2f_lw_axi_master_wvalid,  --                  .wvalid
			h2f_lw_WREADY            => hps_0_h2f_lw_axi_master_wready,  --                  .wready
			h2f_lw_BID               => hps_0_h2f_lw_axi_master_bid,     --                  .bid
			h2f_lw_BRESP             => hps_0_h2f_lw_axi_master_bresp,   --                  .bresp
			h2f_lw_BVALID            => hps_0_h2f_lw_axi_master_bvalid,  --                  .bvalid
			h2f_lw_BREADY            => hps_0_h2f_lw_axi_master_bready,  --                  .bready
			h2f_lw_ARID              => hps_0_h2f_lw_axi_master_arid,    --                  .arid
			h2f_lw_ARADDR            => hps_0_h2f_lw_axi_master_araddr,  --                  .araddr
			h2f_lw_ARLEN             => hps_0_h2f_lw_axi_master_arlen,   --                  .arlen
			h2f_lw_ARSIZE            => hps_0_h2f_lw_axi_master_arsize,  --                  .arsize
			h2f_lw_ARBURST           => hps_0_h2f_lw_axi_master_arburst, --                  .arburst
			h2f_lw_ARLOCK            => hps_0_h2f_lw_axi_master_arlock,  --                  .arlock
			h2f_lw_ARCACHE           => hps_0_h2f_lw_axi_master_arcache, --                  .arcache
			h2f_lw_ARPROT            => hps_0_h2f_lw_axi_master_arprot,  --                  .arprot
			h2f_lw_ARVALID           => hps_0_h2f_lw_axi_master_arvalid, --                  .arvalid
			h2f_lw_ARREADY           => hps_0_h2f_lw_axi_master_arready, --                  .arready
			h2f_lw_RID               => hps_0_h2f_lw_axi_master_rid,     --                  .rid
			h2f_lw_RDATA             => hps_0_h2f_lw_axi_master_rdata,   --                  .rdata
			h2f_lw_RRESP             => hps_0_h2f_lw_axi_master_rresp,   --                  .rresp
			h2f_lw_RLAST             => hps_0_h2f_lw_axi_master_rlast,   --                  .rlast
			h2f_lw_RVALID            => hps_0_h2f_lw_axi_master_rvalid,  --                  .rvalid
			h2f_lw_RREADY            => hps_0_h2f_lw_axi_master_rready   --                  .rready
		);

	sysid_qsys_0 : component soc_system_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component soc_system_mm_interconnect_0
		port map (
			hps_0_h2f_lw_axi_master_awid                                        => hps_0_h2f_lw_axi_master_awid,                                  --                                       hps_0_h2f_lw_axi_master.awid
			hps_0_h2f_lw_axi_master_awaddr                                      => hps_0_h2f_lw_axi_master_awaddr,                                --                                                              .awaddr
			hps_0_h2f_lw_axi_master_awlen                                       => hps_0_h2f_lw_axi_master_awlen,                                 --                                                              .awlen
			hps_0_h2f_lw_axi_master_awsize                                      => hps_0_h2f_lw_axi_master_awsize,                                --                                                              .awsize
			hps_0_h2f_lw_axi_master_awburst                                     => hps_0_h2f_lw_axi_master_awburst,                               --                                                              .awburst
			hps_0_h2f_lw_axi_master_awlock                                      => hps_0_h2f_lw_axi_master_awlock,                                --                                                              .awlock
			hps_0_h2f_lw_axi_master_awcache                                     => hps_0_h2f_lw_axi_master_awcache,                               --                                                              .awcache
			hps_0_h2f_lw_axi_master_awprot                                      => hps_0_h2f_lw_axi_master_awprot,                                --                                                              .awprot
			hps_0_h2f_lw_axi_master_awvalid                                     => hps_0_h2f_lw_axi_master_awvalid,                               --                                                              .awvalid
			hps_0_h2f_lw_axi_master_awready                                     => hps_0_h2f_lw_axi_master_awready,                               --                                                              .awready
			hps_0_h2f_lw_axi_master_wid                                         => hps_0_h2f_lw_axi_master_wid,                                   --                                                              .wid
			hps_0_h2f_lw_axi_master_wdata                                       => hps_0_h2f_lw_axi_master_wdata,                                 --                                                              .wdata
			hps_0_h2f_lw_axi_master_wstrb                                       => hps_0_h2f_lw_axi_master_wstrb,                                 --                                                              .wstrb
			hps_0_h2f_lw_axi_master_wlast                                       => hps_0_h2f_lw_axi_master_wlast,                                 --                                                              .wlast
			hps_0_h2f_lw_axi_master_wvalid                                      => hps_0_h2f_lw_axi_master_wvalid,                                --                                                              .wvalid
			hps_0_h2f_lw_axi_master_wready                                      => hps_0_h2f_lw_axi_master_wready,                                --                                                              .wready
			hps_0_h2f_lw_axi_master_bid                                         => hps_0_h2f_lw_axi_master_bid,                                   --                                                              .bid
			hps_0_h2f_lw_axi_master_bresp                                       => hps_0_h2f_lw_axi_master_bresp,                                 --                                                              .bresp
			hps_0_h2f_lw_axi_master_bvalid                                      => hps_0_h2f_lw_axi_master_bvalid,                                --                                                              .bvalid
			hps_0_h2f_lw_axi_master_bready                                      => hps_0_h2f_lw_axi_master_bready,                                --                                                              .bready
			hps_0_h2f_lw_axi_master_arid                                        => hps_0_h2f_lw_axi_master_arid,                                  --                                                              .arid
			hps_0_h2f_lw_axi_master_araddr                                      => hps_0_h2f_lw_axi_master_araddr,                                --                                                              .araddr
			hps_0_h2f_lw_axi_master_arlen                                       => hps_0_h2f_lw_axi_master_arlen,                                 --                                                              .arlen
			hps_0_h2f_lw_axi_master_arsize                                      => hps_0_h2f_lw_axi_master_arsize,                                --                                                              .arsize
			hps_0_h2f_lw_axi_master_arburst                                     => hps_0_h2f_lw_axi_master_arburst,                               --                                                              .arburst
			hps_0_h2f_lw_axi_master_arlock                                      => hps_0_h2f_lw_axi_master_arlock,                                --                                                              .arlock
			hps_0_h2f_lw_axi_master_arcache                                     => hps_0_h2f_lw_axi_master_arcache,                               --                                                              .arcache
			hps_0_h2f_lw_axi_master_arprot                                      => hps_0_h2f_lw_axi_master_arprot,                                --                                                              .arprot
			hps_0_h2f_lw_axi_master_arvalid                                     => hps_0_h2f_lw_axi_master_arvalid,                               --                                                              .arvalid
			hps_0_h2f_lw_axi_master_arready                                     => hps_0_h2f_lw_axi_master_arready,                               --                                                              .arready
			hps_0_h2f_lw_axi_master_rid                                         => hps_0_h2f_lw_axi_master_rid,                                   --                                                              .rid
			hps_0_h2f_lw_axi_master_rdata                                       => hps_0_h2f_lw_axi_master_rdata,                                 --                                                              .rdata
			hps_0_h2f_lw_axi_master_rresp                                       => hps_0_h2f_lw_axi_master_rresp,                                 --                                                              .rresp
			hps_0_h2f_lw_axi_master_rlast                                       => hps_0_h2f_lw_axi_master_rlast,                                 --                                                              .rlast
			hps_0_h2f_lw_axi_master_rvalid                                      => hps_0_h2f_lw_axi_master_rvalid,                                --                                                              .rvalid
			hps_0_h2f_lw_axi_master_rready                                      => hps_0_h2f_lw_axi_master_rready,                                --                                                              .rready
			clk_0_clk_clk                                                       => clk_clk,                                                       --                                                     clk_0_clk.clk
			Easy_Driver_Y_reset_reset_bridge_in_reset_reset                     => rst_controller_reset_out_reset,                                --                     Easy_Driver_Y_reset_reset_bridge_in_reset.reset
			hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                            -- hps_0_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
			Easy_Driver_X_avalon_slave_dir_write                                => mm_interconnect_0_easy_driver_x_avalon_slave_dir_write,        --                                Easy_Driver_X_avalon_slave_dir.write
			Easy_Driver_X_avalon_slave_dir_read                                 => mm_interconnect_0_easy_driver_x_avalon_slave_dir_read,         --                                                              .read
			Easy_Driver_X_avalon_slave_dir_readdata                             => mm_interconnect_0_easy_driver_x_avalon_slave_dir_readdata,     --                                                              .readdata
			Easy_Driver_X_avalon_slave_dir_writedata                            => mm_interconnect_0_easy_driver_x_avalon_slave_dir_writedata,    --                                                              .writedata
			Easy_Driver_X_avalon_slave_duty_write                               => mm_interconnect_0_easy_driver_x_avalon_slave_duty_write,       --                               Easy_Driver_X_avalon_slave_duty.write
			Easy_Driver_X_avalon_slave_duty_read                                => mm_interconnect_0_easy_driver_x_avalon_slave_duty_read,        --                                                              .read
			Easy_Driver_X_avalon_slave_duty_readdata                            => mm_interconnect_0_easy_driver_x_avalon_slave_duty_readdata,    --                                                              .readdata
			Easy_Driver_X_avalon_slave_duty_writedata                           => mm_interconnect_0_easy_driver_x_avalon_slave_duty_writedata,   --                                                              .writedata
			Easy_Driver_X_avalon_slave_period_write                             => mm_interconnect_0_easy_driver_x_avalon_slave_period_write,     --                             Easy_Driver_X_avalon_slave_period.write
			Easy_Driver_X_avalon_slave_period_read                              => mm_interconnect_0_easy_driver_x_avalon_slave_period_read,      --                                                              .read
			Easy_Driver_X_avalon_slave_period_readdata                          => mm_interconnect_0_easy_driver_x_avalon_slave_period_readdata,  --                                                              .readdata
			Easy_Driver_X_avalon_slave_period_writedata                         => mm_interconnect_0_easy_driver_x_avalon_slave_period_writedata, --                                                              .writedata
			Easy_Driver_X_avalon_slave_step_write                               => mm_interconnect_0_easy_driver_x_avalon_slave_step_write,       --                               Easy_Driver_X_avalon_slave_step.write
			Easy_Driver_X_avalon_slave_step_read                                => mm_interconnect_0_easy_driver_x_avalon_slave_step_read,        --                                                              .read
			Easy_Driver_X_avalon_slave_step_readdata                            => mm_interconnect_0_easy_driver_x_avalon_slave_step_readdata,    --                                                              .readdata
			Easy_Driver_X_avalon_slave_step_writedata                           => mm_interconnect_0_easy_driver_x_avalon_slave_step_writedata,   --                                                              .writedata
			Easy_Driver_Y_avalon_slave_dir_write                                => mm_interconnect_0_easy_driver_y_avalon_slave_dir_write,        --                                Easy_Driver_Y_avalon_slave_dir.write
			Easy_Driver_Y_avalon_slave_dir_read                                 => mm_interconnect_0_easy_driver_y_avalon_slave_dir_read,         --                                                              .read
			Easy_Driver_Y_avalon_slave_dir_readdata                             => mm_interconnect_0_easy_driver_y_avalon_slave_dir_readdata,     --                                                              .readdata
			Easy_Driver_Y_avalon_slave_dir_writedata                            => mm_interconnect_0_easy_driver_y_avalon_slave_dir_writedata,    --                                                              .writedata
			Easy_Driver_Y_avalon_slave_duty_write                               => mm_interconnect_0_easy_driver_y_avalon_slave_duty_write,       --                               Easy_Driver_Y_avalon_slave_duty.write
			Easy_Driver_Y_avalon_slave_duty_read                                => mm_interconnect_0_easy_driver_y_avalon_slave_duty_read,        --                                                              .read
			Easy_Driver_Y_avalon_slave_duty_readdata                            => mm_interconnect_0_easy_driver_y_avalon_slave_duty_readdata,    --                                                              .readdata
			Easy_Driver_Y_avalon_slave_duty_writedata                           => mm_interconnect_0_easy_driver_y_avalon_slave_duty_writedata,   --                                                              .writedata
			Easy_Driver_Y_avalon_slave_period_write                             => mm_interconnect_0_easy_driver_y_avalon_slave_period_write,     --                             Easy_Driver_Y_avalon_slave_period.write
			Easy_Driver_Y_avalon_slave_period_read                              => mm_interconnect_0_easy_driver_y_avalon_slave_period_read,      --                                                              .read
			Easy_Driver_Y_avalon_slave_period_readdata                          => mm_interconnect_0_easy_driver_y_avalon_slave_period_readdata,  --                                                              .readdata
			Easy_Driver_Y_avalon_slave_period_writedata                         => mm_interconnect_0_easy_driver_y_avalon_slave_period_writedata, --                                                              .writedata
			Easy_Driver_Y_avalon_slave_step_write                               => mm_interconnect_0_easy_driver_y_avalon_slave_step_write,       --                               Easy_Driver_Y_avalon_slave_step.write
			Easy_Driver_Y_avalon_slave_step_read                                => mm_interconnect_0_easy_driver_y_avalon_slave_step_read,        --                                                              .read
			Easy_Driver_Y_avalon_slave_step_readdata                            => mm_interconnect_0_easy_driver_y_avalon_slave_step_readdata,    --                                                              .readdata
			Easy_Driver_Y_avalon_slave_step_writedata                           => mm_interconnect_0_easy_driver_y_avalon_slave_step_writedata,   --                                                              .writedata
			sysid_qsys_0_control_slave_address                                  => mm_interconnect_0_sysid_qsys_0_control_slave_address,          --                                    sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                                 => mm_interconnect_0_sysid_qsys_0_control_slave_readdata          --                                                              .readdata
		);

	rst_controller : component soc_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,         -- reset_in0.reset
			reset_in1      => hps_0_h2f_reset_reset_ports_inv, -- reset_in1.reset
			clk            => clk_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,  -- reset_out.reset
			reset_req      => open,                            -- (terminated)
			reset_req_in0  => '0',                             -- (terminated)
			reset_req_in1  => '0',                             -- (terminated)
			reset_in2      => '0',                             -- (terminated)
			reset_req_in2  => '0',                             -- (terminated)
			reset_in3      => '0',                             -- (terminated)
			reset_req_in3  => '0',                             -- (terminated)
			reset_in4      => '0',                             -- (terminated)
			reset_req_in4  => '0',                             -- (terminated)
			reset_in5      => '0',                             -- (terminated)
			reset_req_in5  => '0',                             -- (terminated)
			reset_in6      => '0',                             -- (terminated)
			reset_req_in6  => '0',                             -- (terminated)
			reset_in7      => '0',                             -- (terminated)
			reset_req_in7  => '0',                             -- (terminated)
			reset_in8      => '0',                             -- (terminated)
			reset_req_in8  => '0',                             -- (terminated)
			reset_in9      => '0',                             -- (terminated)
			reset_req_in9  => '0',                             -- (terminated)
			reset_in10     => '0',                             -- (terminated)
			reset_req_in10 => '0',                             -- (terminated)
			reset_in11     => '0',                             -- (terminated)
			reset_req_in11 => '0',                             -- (terminated)
			reset_in12     => '0',                             -- (terminated)
			reset_req_in12 => '0',                             -- (terminated)
			reset_in13     => '0',                             -- (terminated)
			reset_req_in13 => '0',                             -- (terminated)
			reset_in14     => '0',                             -- (terminated)
			reset_req_in14 => '0',                             -- (terminated)
			reset_in15     => '0',                             -- (terminated)
			reset_req_in15 => '0'                              -- (terminated)
		);

	rst_controller_001 : component soc_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => hps_0_h2f_reset_reset_ports_inv,    -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_easy_driver_y_avalon_slave_dir_read_ports_inv <= not mm_interconnect_0_easy_driver_y_avalon_slave_dir_read;

	mm_interconnect_0_easy_driver_y_avalon_slave_dir_write_ports_inv <= not mm_interconnect_0_easy_driver_y_avalon_slave_dir_write;

	mm_interconnect_0_easy_driver_x_avalon_slave_dir_read_ports_inv <= not mm_interconnect_0_easy_driver_x_avalon_slave_dir_read;

	mm_interconnect_0_easy_driver_x_avalon_slave_dir_write_ports_inv <= not mm_interconnect_0_easy_driver_x_avalon_slave_dir_write;

	mm_interconnect_0_easy_driver_y_avalon_slave_duty_read_ports_inv <= not mm_interconnect_0_easy_driver_y_avalon_slave_duty_read;

	mm_interconnect_0_easy_driver_y_avalon_slave_duty_write_ports_inv <= not mm_interconnect_0_easy_driver_y_avalon_slave_duty_write;

	mm_interconnect_0_easy_driver_x_avalon_slave_duty_read_ports_inv <= not mm_interconnect_0_easy_driver_x_avalon_slave_duty_read;

	mm_interconnect_0_easy_driver_x_avalon_slave_duty_write_ports_inv <= not mm_interconnect_0_easy_driver_x_avalon_slave_duty_write;

	mm_interconnect_0_easy_driver_y_avalon_slave_period_read_ports_inv <= not mm_interconnect_0_easy_driver_y_avalon_slave_period_read;

	mm_interconnect_0_easy_driver_y_avalon_slave_period_write_ports_inv <= not mm_interconnect_0_easy_driver_y_avalon_slave_period_write;

	mm_interconnect_0_easy_driver_x_avalon_slave_period_read_ports_inv <= not mm_interconnect_0_easy_driver_x_avalon_slave_period_read;

	mm_interconnect_0_easy_driver_x_avalon_slave_period_write_ports_inv <= not mm_interconnect_0_easy_driver_x_avalon_slave_period_write;

	mm_interconnect_0_easy_driver_y_avalon_slave_step_read_ports_inv <= not mm_interconnect_0_easy_driver_y_avalon_slave_step_read;

	mm_interconnect_0_easy_driver_y_avalon_slave_step_write_ports_inv <= not mm_interconnect_0_easy_driver_y_avalon_slave_step_write;

	mm_interconnect_0_easy_driver_x_avalon_slave_step_read_ports_inv <= not mm_interconnect_0_easy_driver_x_avalon_slave_step_read;

	mm_interconnect_0_easy_driver_x_avalon_slave_step_write_ports_inv <= not mm_interconnect_0_easy_driver_x_avalon_slave_step_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	hps_0_h2f_reset_reset_ports_inv <= not hps_0_h2f_reset_reset;

end architecture rtl; -- of soc_system
